
entity 